package constantsMIDI;
    parameter NOTE_ON = 1;
    parameter NOTE_OFF = 0;
endpackage